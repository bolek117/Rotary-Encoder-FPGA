//-----------------------------------------------------------------------------
//
// Title       : rotaryQueue_tb
// Design      : project2
// Author      : 
// Company     : 
//
//-----------------------------------------------------------------------------
//
// File        : D:\Program Files (x86)\Aldec\Designs\proj2\project2\src\rotaryQueue_tb.v
// Generated   : Wed Feb 12 18:15:47 2014
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {rotaryQueue_tb}}
module rotaryQueue_tb;

	

endmodule
